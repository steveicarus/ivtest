// Copyright (c) 2006 Stephen Williams
//
//    This source code is free software; you can redistribute it
//    and/or modify it in source code form under the terms of the GNU
//    General Public License as published by the Free Software
//    Foundation; either version 2 of the License, or (at your option)
//    any later version.
//
//    This program is distributed in the hope that it will be useful,
//    but WITHOUT ANY WARRANTY; without even the implied warranty of
//    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
//    GNU General Public License for more details.
//
//    You should have received a copy of the GNU General Public License
//    along with this program; if not, write to the Free Software
//    Foundation, Inc., 59 Temple Place - Suite 330, Boston, MA 02111-1307, USA
//

module main;

   reg [7:0] mem [0:1];

   initial begin
      mem[0] = 0;
      mem[1] = 1;
      $memmonitor(mem);

      #1 mem[0] = 4;
      #1 mem[1] = 5;
      #1 $finish;
   end

endmodule // main
