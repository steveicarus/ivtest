`timescale 1ns/1ps
module top;
`timescale 1us/1ns
endmodule


