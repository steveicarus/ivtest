module top;
  int bound = 2;
  string q_str1 [$:-1];
  string q_str2 [$:bound];

  initial $display("FAILED");
endmodule : top
