module tb;
initial $finish;
final $display("In final statement.");
endmodule
