module tb;
final $display("In final statement.");
endmodule
