module top;

  initial begin
    $display("Output a slash \\.");
    $display("Output a double slash \\\\.");
  end
endmodule

 	  	 
