module top;
  int bound = 2;
  int q_vec1 [$:-1];
  int q_vec2 [$:bound];

  initial $display("FAILED");
endmodule : top
