module top;
  initial begin
    $display("PASSED");
  end;
endmodule
