// Copyright (c) 2015 CERN
// Maciej Suminski <maciej.suminski@cern.ch>
//
// This source code is free software; you can redistribute it
// and/or modify it in source code form under the terms of the GNU
// General Public License as published by the Free Software
// Foundation; either version 2 of the License, or (at your option)
// any later version.
//
// This program is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
// GNU General Public License for more details.
//
// You should have received a copy of the GNU General Public License
// along with this program; if not, write to the Free Software
// Foundation, Inc., 59 Temple Place - Suite 330, Boston, MA 02111-1307, USA


// Test for constant arrays access

module constant_array_test;
reg logic [7:0] out_word;
reg logic [2:0] index;
constant_array dut(index, out_word);

initial begin
  index = 2;
  #1;       // wait for signal assignments

  if(out_word !== 16)
  begin
    $display("FAILED 1");
    $finish();
  end

  index = 4;
  #1;

  if(out_word !== 64)
  begin
    $display("FAILED 2");
    $finish();
  end

  if(dut.test_a !== 32)
  begin
    $display("FAILED 3");
    $finish();
  end

  if(dut.test_b !== 4)
  begin
    $display("FAILED 4");
    $finish();
  end

  if(dut.test_c !== 3'b100)
  begin
    $display("FAILED 5");
    $finish();
  end

  if(dut.test_d !== 1'b1)
  begin
    $display("FAILED 6");
    $finish();
  end

  $display("PASSED");
end
endmodule
