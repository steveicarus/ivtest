module top();

  register loop();
  process signal();
  
endmodule // top

module register();

endmodule // register

module process();

  initial $display("PASSED");
  
endmodule // process
