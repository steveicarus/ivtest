//---------------------------------------------------------------------------
// 
//---------------------------------------------------------------------------
 module xor_try;

   (* ivl_do_not_elide *) reg unused;
   initial $sn;
 endmodule

