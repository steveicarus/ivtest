module testbench;
foo #(ASDF) bar(); 
endmodule

module foo #(parameter A=1);
endmodule
