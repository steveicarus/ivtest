
module sub8(output wire [7:0] out, input wire [7:0] A, input wire [7:0] B);

   assign out = A - B;

endmodule
